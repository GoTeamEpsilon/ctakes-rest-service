// CUI|TUI|Text|preferredTerm
// CUI|TUI|Text|preferredTerm
C0201838|T059|Albumin measurement
C0202202|T059|Protein measurement
C0201850|T059|Alkaline phosphatase measurement
C0201836|T059|Alanine aminotransferase measurement
C0201836|T059|ALT
C0201899|T059|AST
C0201899|T059|Aspartate aminotransferase measurement
C0201913|T059|Bilirubin, total measurement|bilirubin
C0036808|T059|Serum Indirect (Unconjugated) Bilirubin Test
C0858048|T059|Bilirubin, Direct
C0201973|T059|Total CK
C0201973|T059|Creatine kinase measurement
C0523584|T059|CK-MB
C0523584|T059|Creatine kinase MB measurement
C0523584|T059|CKMB
C0523584|T059|Creatine kinase MB measurement
C0023508|T059|White Blood Cell Count procedure
C0023508|T059|white count
C0201803|T059|Osmolality Measurement
C0201803|T059|osmolality
C0017654|T060|Glomerular Filtration Rate
C0017654|T060|GFR
C0588466|T059|Red blood cells urine (lab test)
C0588466|T059|RBC, UA
C0023508|T059|White Blood Cell Count procedure
C0919738|T059|White blood cells urine (lab test)
C0919738|T059|WBC, UA
C0201837|T059|Albumin/Globulin ratio
C0201837|T059|A/G Ratio
C0373670|T059|Lipase measurement
C0373670|T059|Lipase
C0033707|T059|Protime
C0033707|T059|Prothrombin time assay
C0525032|T059|International Normalized Ratio
C0525032|T059|INR
C1443182|T059|Calculated (procedure)
C1443182|T059|Calc
C0337443|T059|Na
C0337443|T059|sodium
C0337443|T059|Sodium measurement
C0202194|T059|potassium
C0202194|T059|Potassium measurement
C0202194|T059|pot
C0202194|T059|pota
C0202194|T059|potas
C0003074|T201|Anion Gap
C0202230|T059|TSH
C0202230|T059|Thyroid stimulating hormone measurement
C1171408|T059|High density/low density lipoprotein ratio measurement
C1171408|T059|LDL/HDL
C0518015|T059|hemoglobin
C0518015|T059|Hemoglobin measurement
C0032181|T059|platelet count
C0032181|T059|Platelet Count measurement
C0018935|T059|Hematocrit procedure
C0018935|T059|hematocrit
C0201657|T059|CRP
C0201657|T059|C-reactive protein measurement
C1535922|T059|procalcitonin
C1535922|T059|Procalcitonin measurement
C0202115|T059|lactate
C0202115|T059|Lactic acid measurement
C0202225|T059|T4 free measurement
C0202225|T059|free T4
C0201934|T059|Cardiac enzymes measurement
C0201934|T059|cardiac enzymes
C0337438|T059|glucose
C0337438|T059|Glucose measurement
C0201802|T059|specific gravity
C0200635|T059|Lymphocyte Count measurement
C0201802|T059|Specific gravity measurement
C0200635|T059|lymphocytes
C0005845|T059|Blood urea nitrogen measurement
C0005845|T059|BUN
C0201975|T059|Creatinine measurement
C0201975|T059|creatinine
C1305866|T060|weight
C1305866|T060|Weighing patient
C1305855|T201|BMI
C1305855|T201|Body mass index
C0489786|T032|Height
C0489786|T032|Ht
C0302353|T059|Serum potassium measurement
C0302353|T059|Serum potassium
C0523891|T059|Serum sodium measurement
C0523891|T059|Serum sodium
C0600061|T033|Serum creatinine level
C0600061|T033|SERUM CREATININE
C0728876|T059|Serum calcium measurement
C0728876|T059|Serum calcium
C0202178|T059|Phosphorus measurement
C0202178|T059|Phosphorus Test
C0041942|T109|Urea
C0523465|T059|SERUM ALBUMIN measurement
C0523465|T059|SERUM ALBUMIN 
C0201916|T059|DIRECT BILIRUBIN 
C0201916|T059|Bilirubin, direct measurement
C0428326|T059|SGPT - blood measurement  
C0428326|T059|SGPT
C0201913|T059|BILIRUBIN
C0201913|T059|Bilirubin, total measurement
C0151415|T033|SGOT
C0151415|T033|SGOT,patient value
C0555903|T059|TOTAL PROTEIN
C0555903|T059|Total protein measurement
C0201850|T059|ALKALINE PHOSPHATASE
C0201850|T059|ALKALINE PHOSPHATASE measurement
C2677004|T033|Increased serum gamma-GGT
C2677004|T033|SERUM GGT
C0033706|T123|Prothrombin
C0150012|T033|Does Patient Have A Difficult Airway/Aspiration Risk?
C0150012|T033|At risk for aspiration
C0553700|T033|Actual blood loss
C0282638|T061|Antibiotic Prophylaxis
C0282638|T061|Has antibiotic prophylaxis been given within the last 60 minutes?
C0853245|T061|Has DVT prophylaxis been administered
C0853245|T061|DVT prophylaxis
C0201617|T059|PLT
C0201617|T059|Primed lymphocyte test
C4055231|T185|maxCD
C4055231|T185|newCD
C3248554|T201|post-operative day 1
C3248554|T201|post-operative day 2
C3248554|T201|post-operative day 3
C3248554|T201|post-operative day 4
C3248554|T201|post-operative day 5
C3248554|T201|post-operative day 6
C3248554|T201|post-operative day 7
C3248554|T201|post operative day 1
C3248554|T201|post operative day 3
C3248554|T201|post operative day 4
C3248554|T201|post operative day 5
C3248554|T201|post operative day 6
C3248554|T201|post operative day 7
C3248554|T201|pod 1
C3248554|T201|pod 2
C3248554|T201|pod 3
C3248554|T201|pod 4
C3248554|T201|pod 5
C3248554|T201|pod 6
C3248554|T201|pod 7
C3248554|T201|POD 1
C3248554|T201|POD 2
C3248554|T201|POD 3
C3248554|T201|POD 4
C3248554|T201|POD 5
C3248554|T201|POD 6
C3248554|T201|POD 7
C3248561|T201|post-operative day 8
C3248561|T201|post-operative day 9
C3248561|T201|post-operative day 10
C3248561|T201|post-operative day 11
C3248561|T201|post-operative day 12
C3248561|T201|post-operative day 13
C3248561|T201|post-operative day 14
C3248561|T201|post operative day 8
C3248561|T201|post operative day 9
C3248561|T201|post operative day 10
C3248561|T201|post operative day 11
C3248561|T201|post operative day 12
C3248561|T201|post operative day 13
C3248561|T201|post operative day 14
C3248561|T201|pod 8
C3248561|T201|pod 9
C3248561|T201|pod 10
C3248561|T201|pod 11
C3248561|T201|pod 12
C3248561|T201|pod 13
C3248561|T201|pod 14
C3248561|T201|POD 8
C3248561|T201|POD 9
C3248561|T201|POD 10
C3248561|T201|POD 11
C3248561|T201|POD 12
C3248561|T201|POD 13
C3248561|T201|POD 14
C0871470|T201|Blood Pressure
C0871470|T201|Systolic Blood Pressure
C0871470|T201|Sys Blood Pressure
C0871470|T201|SBP
C0871470|T201|Sys BP
C0428883|T201|Diastolic Blood Pressure
C0428883|T201|Dia Blood Pressure
C0428883|T201|DBP
C0428883|T201|Dia BP
C0429774|T201|Residual urine volume
C0429774|T201|Residual urine vol
C0429774|T201|urine volume
C0429774|T201|urine vol
C0429774|T201|Res urine volume
C0429774|T201|Res urine vol
C0041657|T201|Unconscious State
C0041657|T201|Unconscious
C0426498|T201|Dry tongue
C0234421|T201|Conscious
C0005903|T201|Temperature
C0005903|T201|Temp
C1321898|T201|Blood in stool
C1321898|T201|Blood stool



	

































 












